----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 02/10/2017 11:07:04 AM
-- Design Name: 
-- Module Name: Video_Box - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity image_overlay is
port (
    --reg in
     slv_reg0 : in std_logic_vector(31 downto 0);  -- x
     slv_reg1 : in std_logic_vector(31 downto 0);  -- y
     slv_reg2 : in std_logic_vector(31 downto 0);  -- width
     slv_reg3 : in std_logic_vector(31 downto 0);  -- height
     slv_reg4 : in std_logic_vector(31 downto 0);
     slv_reg5 : in std_logic_vector(31 downto 0);  
     slv_reg6 : in std_logic_vector(31 downto 0);  
     slv_reg7 : in std_logic_vector(31 downto 0);    
     
    --reg out
    slv_reg0out : out std_logic_vector(31 downto 0);  
    slv_reg1out : out std_logic_vector(31 downto 0);  
    slv_reg2out : out std_logic_vector(31 downto 0);  
    slv_reg3out : out std_logic_vector(31 downto 0);  
    slv_reg4out : out std_logic_vector(31 downto 0);
    slv_reg5out : out std_logic_vector(31 downto 0);  
    slv_reg6out : out std_logic_vector(31 downto 0);  
    slv_reg7out : out std_logic_vector(31 downto 0);
    
    --Bus Clock
    CLK : in std_logic;
    --Video
    RGB_IN_I : in std_logic_vector(23 downto 0); -- Parallel video data (required)
    VDE_IN_I : in std_logic; -- Active video Flag (optional)
    HB_IN_I : in std_logic; -- Horizontal blanking signal (optional)
    VB_IN_I : in std_logic; -- Vertical blanking signal (optional)
    HS_IN_I : in std_logic; -- Horizontal sync signal (optional)
    VS_IN_I : in std_logic; -- Veritcal sync signal (optional)
    ID_IN_I : in std_logic; -- Field ID (optional)
    --  additional ports here
    RGB_IN_O : out std_logic_vector(23 downto 0); -- Parallel video data (required)
    VDE_IN_O : out std_logic; -- Active video Flag (optional)
    HB_IN_O : out std_logic; -- Horizontal blanking signal (optional)
    VB_IN_O : out std_logic; -- Vertical blanking signal (optional)
    HS_IN_O : out std_logic; -- Horizontal sync signal (optional)
    VS_IN_O : out std_logic; -- Veritcal sync signal (optional)
    ID_IN_O : out std_logic; -- Field ID (optional)
    
    PIXEL_CLK_IN : in std_logic;
    
    X_Cord : in std_logic_vector(15 downto 0);
    Y_Cord : in std_logic_vector(15 downto 0)

);
end image_overlay;

architecture Behavioral of image_overlay is


--signal red, blue, green : std_logic_vector(7 downto 0);
--signal lred, lblue, lgreen : std_logic_vector(7 downto 0);
	
signal rgb_next : std_logic_vector(23 downto 0);
signal use_image : std_logic;
signal image_next_index : integer := 0;
signal image_next_pixel : std_logic_vector(23 downto 0);

signal int_X_Coord : unsigned(15 downto 0);
signal int_Y_Coord : unsigned(15 downto 0);
signal int_X_Orig : unsigned(31 downto 0);
signal int_Y_Orig : unsigned(31 downto 0);
signal img_width : unsigned(31 downto 0);
signal img_height : unsigned(31 downto 0);

constant N : integer := 14;
type ram_type is array(0 to 2**N-1) of std_logic_vector(23 downto 0);

signal image : ram_type := (
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FEFBFF", x"FCFAFF", x"FFFFFC", x"FFFFF9", x"FEFFFF", x"F9FEFF", x"FEFFFC", x"FFFFF1", x"FFFCFF", x"FEFDFA", x"FFFEFF", x"FFF8FF", x"FBFFFC", x"FEFEFE", x"FFFEFB", x"FFFEF9", x"EFF2F9", x"E7EBF1", x"E9ECF2", x"F6FAFF", x"FFFFFC", x"FFFCFE", x"FEFFFC", x"F8FEF6", x"FFFEFF", x"FCFDFA", x"FEFEFE", x"FCFBFF", x"FCFDFA", x"F9FEFF", x"FDFFFB", x"FDFEF6", x"FEFDF7", x"FFFCFF", x"FFFEFF", x"FFFCFE", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FEFFFC", x"FEFFFF", x"FCFCFC", x"FEFEFF", x"FFFFF9", x"FAFFF5", x"FEFCFF", x"FFF8FF", x"F7F7FF", x"868AAF", x"26385D", x"0E2843", x"1D2F55", x"43577A", x"697E95", x"8FA2B3", x"BABFC7", x"CAD0D7", x"C4CAD1", x"AEB4BB", x"8195A7", x"576B8A", x"2F416A", x"15244B", x"1A3353", x"475377", x"C2C5DC", x"FDFFFE", x"FFFCFF", x"F3F8F6", x"FDFFF0", x"FFFEFC", x"FFFFFF", x"FDFFFE", x"FDFFFB", x"FDFFFB", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFDF9", x"FFFEFF", x"FFFEFF", x"FEFFF2", x"FBFFFC", x"9399B3", x"1B2450", x"1F3158", x"9BA3BB", x"FEFBFC", x"FEFFF9", x"FAFFFF", x"FFFCFB", x"FEFCFF", x"FEFFFF", x"FBFAFF", x"FDFEFF", x"FEFFFF", x"FEFFFF", x"FDFEFF", x"FEFCFF", x"FEFFFF", x"FEFBFC", x"FFFAF6", x"F0F5F6", x"FFFEF7", x"EEF2FE", x"606A88", x"122043", x"3B4269", x"E5E7F6", x"FCFCFF", x"FEFFF7", x"FFFEFF", x"FFFCFE", x"FFFDF4", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"F7F3FC", x"FBFFFA", x"B5C0CF", x"171C3D", x"455473", x"F5FBFF", x"FFFFF5", x"FEFFEE", x"FAFFFF", x"F5FDFA", x"B9C4D0", x"5C6986", x"22355C", x"081439", x"010930", x"06032C", x"000029", x"01002A", x"000029", x"01002A", x"01042B", x"061037", x"0E1C42", x"3B5079", x"838FA8", x"E4EEF0", x"F6FEFB", x"F4FDFF", x"FBFAF4", x"FFFFFA", x"B2C1CB", x"13203E", x"454C6A", x"F1FDFB", x"FDFFFB", x"FFFBFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FEFBFF", x"F7F9F2", x"FEFFF9", x"FEFEFB", x"FEFCFF", x"FFFFFA", x"FAFFF9", x"FFFBFF", x"5F6A84", x"161C41", x"E3EAEA", x"FFFEFF", x"FFFFFC", x"FFFEFA", x"ADB2CB", x"28325D", x"00072D", x"010E33", x"061941", x"07214A", x"021D47", x"021A48", x"042046", x"011C48", x"021E48", x"021E43", x"071E49", x"031B49", x"021D45", x"071E45", x"031E44", x"022041", x"011B41", x"001039", x"00002D", x"070D38", x"575F86", x"E9E8EB", x"FFFFF5", x"FAFBFF", x"F5FEF5", x"6D7189", x"151C42", x"D6ECF1", x"FFFFFF", x"FEFFF2", x"FFFCFF", x"FFFEFF", x"FDFFF7", x"FEFFFC", x"FFFFFF", x"FFFCFE", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFC", x"FFFCFF", x"FEFBFF", x"FFFEFF", x"FAFBF5", x"FCFAFB", x"58667E", x"272C4D", x"F9FCFF", x"F6FDFF", x"FAFDF6", x"BCB3C9", x"192240", x"000235", x"081648", x"022040", x"061D46", x"011B43", x"011840", x"091B48", x"0A1E48", x"031942", x"021F46", x"021D41", x"071E49", x"081F40", x"051C4A", x"021F3B", x"021E43", x"031E44", x"061F48", x"011943", x"021F44", x"011B45", x"021F42", x"021E3F", x"08214A", x"050D40", x"000028", x"4B5D77", x"FFFEFF", x"FBFCFF", x"FAFFFF", x"B0B1C7", x"0C1735", x"EEF5F5", x"F6FBFA", x"FFFBFF", x"FFFCFF", x"FBFAF7", x"FFFEFF", x"FEFFF7", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFC", x"FFFEFF", x"FCFDFA", x"F8FEF6", x"A4AFBB", x"131B42", x"F6F9F5", x"FEFFF9", x"FBFDF5", x"646E91", x"000728", x"051945", x"061B44", x"081E42", x"031D41", x"021B44", x"081F48", x"071E45", x"092046", x"021D43", x"000E32", x"011436", x"021F4C", x"132E52", x"020F38", x"071D4B", x"021D44", x"0F1D47", x"0C193E", x"011B45", x"021D3F", x"051C42", x"071941", x"0A1947", x"011B46", x"0A1C4A", x"092046", x"041C43", x"021B41", x"091D44", x"010930", x"0E1D40", x"DAD7E5", x"FFFFFA", x"FFFFFA", x"9CA6B7", x"131A3C", x"F5FFFF", x"FBFEFC", x"FFFEFF", x"FFFFF1", x"F7F7FF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"F6F6F4", x"F7F7F7", x"F0F7FF", x"0B1224", x"DBDFED", x"F7F6FC", x"FAFFFF", x"666B87", x"000229", x"021F4B", x"0A1E42", x"011B46", x"041F47", x"011A44", x"081E4A", x"011942", x"011B3A", x"011332", x"283E68", x"01163C", x"929BBF", x"3A4663", x"061C4A", x"05102C", x"EEFBFF", x"090927", x"0F2048", x"2A3D62", x"384660", x"081A49", x"000D2D", x"575E88", x"727FA7", x"607091", x"000C28", x"022049", x"011B45", x"041F44", x"021D45", x"011A49", x"041D40", x"021E48", x"04103C", x"031232", x"DADDF5", x"FBFFFF", x"FFFCFF", x"2F4158", x"798295", x"FEFFFF", x"FFFCFF", x"FDFFF0", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FEFFFA", x"F8FFFF", x"FEF7FF", x"FEFFF7", x"FFFCFF", x"97A6B3", x"333561", x"FFFFEE", x"FEFDF6", x"A49FC2", x"00062C", x"03204A", x"0A1E4A", x"091D3D", x"021950", x"041F3A", x"0B0D44", x"020927", x"061444", x"022145", x"181340", x"FFFEEF", x"000026", x"061E41", x"000626", x"4E5672", x"04214A", x"000E39", x"647996", x"F9FEFF", x"040126", x"112C4C", x"1D2F52", x"071941", x"D5E5F0", x"05002D", x"01153F", x"00001A", x"D1D6E1", x"0A1B4D", x"041D42", x"021E43", x"022047", x"031A51", x"021F4A", x"071B3B", x"021F4C", x"031C42", x"06113D", x"182143", x"F5FDFF", x"FFFDF1", x"FFFBFF", x"000D2A", x"FEFFFF", x"FFFEF7", x"FAFFFE", x"FFFEFC", x"F9FFFE", x"FFFBFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FEFEF1", x"FEFEFF", x"FEFBFC", x"F6FFF7", x"18244A", x"D6D4E8", x"F6FEFB", x"FBF7FF", x"10112F", x"071D40", x"0A1E48", x"061D44", x"071C43", x"021D41", x"021D43", x"000C30", x"9F9FBA", x"B8BABE", x"FFF3FC", x"080026", x"091C3F", x"BBC0D7", x"0A1A4C", x"04214A", x"060434", x"8497A3", x"0A1E45", x"0A0735", x"91A7B1", x"000023", x"FFF7FA", x"000430", x"1D3657", x"050A32", x"F6FFFF", x"05153A", x"011C47", x"001241", x"022245", x"021F41", x"011B42", x"041E49", x"01133B", x"627090", x"00022A", x"011A40", x"0A1F4A", x"0C1E3F", x"051A41", x"032048", x"000027", x"7581A9", x"FBFFFF", x"FEFEFF", x"162043", x"DBDDEC", x"FFF8FF", x"F8FCF2", x"FFFDF6", x"F4FFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FCFAFF", x"FFFEFB", x"F4FBFB", x"000025", x"FFFCFF", x"F9F9EF", x"9FA8C3", x"000123", x"031C42", x"011C49", x"021C45", x"021D43", x"04123B", x"022247", x"00072C", x"ADB9D1", x"070B37", x"0A1E45", x"000C29", x"FFFAF6", x"00103D", x"465972", x"3D566E", x"0A204A", x"0B153F", x"9BA3B3", x"071A3F", x"00022A", x"8A9DAD", x"09164A", x"000026", x"F6FFFF", x"061141", x"00002A", x"FFFBF9", x"0A0F36", x"0F1B43", x"BFC8D4", x"5E6F96", x"03153D", x"041E49", x"051B49", x"091439", x"D6DBDC", x"657185", x"05163E", x"010F3A", x"031A48", x"031C45", x"09214E", x"011C47", x"091D45", x"070F37", x"FAF9F2", x"FFFCFB", x"8187A7", x"6B7490", x"F9FFFA", x"FFFBFC", x"FFFDF4", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"F9FAFF", x"F6FFFF", x"090B2F", x"FBFEFA", x"FFFEFF", x"33415E", x"091340", x"081F46", x"021D40", x"0A1E46", x"051C43", x"0F1D47", x"B8B7C8", x"01153C", x"081336", x"727B8E", x"072140", x"021D4B", x"011843", x"FCFBFF", x"000028", x"00052A", x"FFFCFF", x"2B2D4D", x"747591", x"212D4D", x"041E49", x"354571", x"61768C", x"0A1E49", x"0A204A", x"010D36", x"162D4A", x"0C2150", x"51637F", x"656D91", x"000025", x"F1FAFF", x"090021", x"022046", x"021D41", x"091D45", x"0F102D", x"E0EEFE", x"011638", x"021D4B", x"43566B", x"6A7E98", x"02183E", x"011B40", x"061D44", x"091F45", x"072248", x"000029", x"DAE8F7", x"FCFBF6", x"DEEAF6", x"2A3554", x"FFFFFF", x"FEFEFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFF9", x"FFFEFF", x"FFF8FE", x"FAFFF7", x"FFFCFF", x"0C2144", x"FFFFEB", x"FDFEFF", x"060D2E", x"0B1F48", x"051B47", x"021E45", x"031D48", x"000C32", x"172A57", x"000636", x"6F7CA4", x"091D40", x"04002E", x"FAFFF9", x"000A27", x"02214C", x"001034", x"B5C6DD", x"061B41", x"0C2048", x"00042F", x"0A264B", x"000E33", x"051C43", x"011B46", x"061D4A", x"051B45", x"061C46", x"051B45", x"061C46", x"031B49", x"021F45", x"051940", x"020A33", x"3A5782", x"0D1B44", x"081C44", x"022045", x"051C42", x"011A42", x"EDEDED", x"040D45", x"0A1E3D", x"021F40", x"ADC1CA", x"020027", x"011645", x"192B47", x"021B46", x"051C4A", x"031F49", x"041D40", x"000C32", x"9295BE", x"FAF7FB", x"FAFFFF", x"121F3F", x"FEFFF5", x"FEFFFF", x"FFFBF4", x"F2FFFF", x"FFF7FF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"F9FEFC", x"FDFDF2", x"FFFCFF", x"F5FFFF", x"122641", x"FFFEFB", x"FBFFFF", x"000526", x"0E1F46", x"01183F", x"031C47", x"021C42", x"0A1439", x"C7C5D6", x"FFFCFF", x"0B0F2F", x"565D89", x"02204B", x"0C1F47", x"435170", x"FCF7FF", x"595A74", x"A9ACD4", x"060123", x"091F49", x"021C44", x"031B44", x"031F47", x"091B43", x"031A3E", x"091D40", x"091D3D", x"021E46", x"021C44", x"021D45", x"021E46", x"021B3C", x"0A1D43", x"091B42", x"061B42", x"081B43", x"071E45", x"011B43", x"0A1D48", x"061C4A", x"051745", x"FFFBFF", x"000022", x"081C4E", x"000B26", x"39567A", x"02204A", x"071F4E", x"848CB3", x"10243D", x"051C4A", x"021B41", x"031D48", x"062046", x"03143F", x"546E80", x"FBFCFF", x"FFF8FF", x"102043", x"FFFEFC", x"FFFEFF", x"FFF9F6", x"F3FFF6", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FEF7FC", x"FFFEFF", x"F4FFFF", x"0D1438", x"F1FDFB", x"FFFCFE", x"09002E", x"021D41", x"011B45", x"041E49", x"08214A", x"041C43", x"021C3E", x"05143D", x"00092A", x"8C9ABA", x"A0ACC9", x"02183C", x"0E1C4B", x"0A1E4F", x"00002D", x"010C2B", x"071035", x"091A4A", x"021D47", x"061C46", x"021E45", x"021D43", x"021E46", x"021B44", x"061D46", x"031D48", x"031C45", x"011A42", x"021B44", x"031C45", x"071E49", x"011C43", x"061F48", x"021D45", x"011B41", x"061F48", x"011B42", x"032045", x"021F42", x"021E46", x"040326", x"D6E3FF", x"424261", x"CED1FF", x"010C32", x"041E49", x"00002E", x"C0D5DA", x"3B4D68", x"031E46", x"01173A", x"081B48", x"021E3E", x"051B49", x"01183E", x"505E78", x"FFFEFF", x"F8FFFF", x"253054", x"FEFFF6", x"F9FFF6", x"FFFBFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FEFFF7", x"FBFFFF", x"000021", x"FAFFFE", x"FFFAF6", x"000026", x"082050", x"081B4B", x"071E47", x"051A43", x"031F47", x"011B43", x"0A1D44", x"0B1B44", x"051947", x"011439", x"CEDFE0", x"434D69", x"0D1B4A", x"061E41", x"0A204A", x"071E47", x"0A2149", x"032044", x"071B45", x"021C42", x"0B1B44", x"000D35", x"00012E", x"0A183D", x"253D60", x"52688C", x"7A89A3", x"8595AF", x"8190AB", x"72819B", x"3C5075", x"172B4F", x"020D35", x"04002F", x"09183E", x"061A40", x"061D44", x"061F48", x"021D4A", x"021F47", x"032145", x"000E2E", x"01132A", x"020E32", x"0B1540", x"000025", x"EAEBED", x"0C1440", x"8299B4", x"0A2047", x"92A2BD", x"1A2648", x"091F45", x"041E49", x"011946", x"011B3A", x"576B88", x"FBFBF9", x"DFF0F4", x"727A9F", x"FFFCFF", x"F6FDF4", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"F6F9F7", x"FAFEF5", x"FCFBF9", x"FBFFFF", x"F3FEF7", x"000830", x"FAFFFC", x"FFFFFA", x"000827", x"071D44", x"061F48", x"021E4A", x"001344", x"374B72", x"011C47", x"022145", x"071D41", x"041D42", x"051C4B", x"021C40", x"60708C", x"091032", x"011C47", x"0A1E45", x"071D44", x"031940", x"061C48", x"091C49", x"00002E", x"0E1B43", x"8092A6", x"FBFFFF", x"FEFEFB", x"FFFEFF", x"FFFCFF", x"FFFCFB", x"FCFCFF", x"FFFFFF", x"FCFCFF", x"FFFFFF", x"FFFEFF", x"FFFBFF", x"FEFEFF", x"FFFFFA", x"CCD6DF", x"415575", x"000A32", x"0D0E38", x"021A4A", x"051A43", x"081C40", x"062043", x"032045", x"0A1F47", x"172543", x"FEFCFF", x"00081E", x"000732", x"DFD7DC", x"000020", x"9BAEBA", x"09123B", x"021D46", x"071F40", x"041F44", x"021F48", x"05113D", x"91A2C1", x"FFFFF5", x"8495B3", x"E3DDE2", x"FAFBFE", x"F8FCF2", x"FFFCFF", x"FBFFF6", x"FFFEFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FEFFFC", x"FEFEFE", x"FFFAFB", x"F6FEEF", x"475780", x"FFFFFC", x"FFF4F2", x"141C41", x"121E4D", x"011B48", x"022044", x"022244", x"5C7087", x"8693A5", x"000F37", x"022046", x"08204B", x"032045", x"011C47", x"091F46", x"01163F", x"071948", x"021D44", x"0C1A4D", x"081E45", x"021D3D", x"000033", x"787995", x"FBFFFF", x"FFFCFF", x"F8F9EF", x"D4DEE1", x"556384", x"1F2D5C", x"13244F", x"233D5D", x"42557B", x"4E6289", x"4A5E85", x"3A4C72", x"1A3156", x"14224F", x"2C3960", x"8C9CB7", x"FAFFFE", x"FFFEF7", x"FFFEFF", x"DFE5EA", x"202A4B", x"000630", x"0A2048", x"061C48", x"021F44", x"061C46", x"051C4A", x"000F36", x"0D1F45", x"000139", x"F8EAF2", x"DAEBF6", x"000E2C", x"011B4A", x"0F1C45", x"0B1D3F", x"051A43", x"021C42", x"021D41", x"00093A", x"D9E8FF", x"F9FFF7", x"12214D", x"FFFCFE", x"FFFEFF", x"FFFFF0", x"F5F6FB", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FEFFFF", x"FEFBFC", x"FFFEF9", x"EAF3FF", x"8392AD", x"FDFEF7", x"5D7493", x"0A1B44", x"021D42", x"021D47", x"0B1F48", x"031B49", x"01053D", x"A7AFBB", x"C2D8DA", x"02002B", x"02173F", x"011A41", x"021C42", x"011840", x"082148", x"062147", x"041F44", x"0A204A", x"00002D", x"8F9EAD", x"FEFEF1", x"FEFFF5", x"D0DBE4", x"172451", x"2E3963", x"C9CECF", x"FFFBFF", x"FFFCFF", x"FDFEFF", x"FBFEFA", x"FFFCFE", x"FFFEFF", x"FFFCFE", x"FEFBFC", x"FAFFFB", x"FFFEFF", x"FEFBFF", x"FCF7F6", x"767E95", x"0D1649", x"566487", x"F9FBF5", x"F6FFFA", x"FFFEFB", x"2F3261", x"090D35", x"0A1E49", x"021E42", x"031D40", x"021F44", x"071D4A", x"00052E", x"FFFAFF", x"000124", x"071D49", x"021E3C", x"3F4D5C", x"FAFFFF", x"111C40", x"021E48", x"011B40", x"061E4B", x"01002A", x"FFFFFC", x"FFFEF7", x"00022A", x"FBFFFF", x"FFFEFC", x"F8FAF4", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FDFEF7", x"FAFFFF", x"000C26", x"FAFFFF", x"EFEEFB", x"05092E", x"021E45", x"011B3F", x"0C1F47", x"00092A", x"021137", x"091B4D", x"A49FC4", x"212C48", x"FFFBFF", x"667496", x"001039", x"092249", x"031E44", x"011C49", x"071D47", x"000533", x"515E72", x"FEFFFF", x"FEFFFA", x"9295B3", x"111A32", x"CACCDC", x"FEFFF9", x"FCFCFC", x"FFFEF9", x"FFFBFF", x"FFFAFC", x"FFFEFF", x"FEFBFF", x"FFFEFF", x"FFFEFF", x"FFFCFF", x"FFFEFF", x"FFFCFF", x"FFFBFC", x"FFFCFF", x"FFFAFF", x"FCFDFA", x"F9FBF7", x"FBFFFF", x"5C5B78", x"1E2A44", x"FBF8FF", x"FFFEFB", x"EFF6F6", x"070B28", x"091C49", x"0A1E49", x"011B46", x"071C54", x"021E3D", x"051537", x"0A1A40", x"0A1647", x"48657B", x"DEEAF6", x"000029", x"03163A", x"01163B", x"051B45", x"021D40", x"041F47", x"01112D", x"FDFEFF", x"F6FDFF", x"738190", x"FFFFFF", x"FFFFFF", x"FFFFF9", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"F0FFFC", x"FBFEFC", x"364970", x"FFFFFA", x"FFFCFF", x"000327", x"071D43", x"021D4B", x"091A4A", x"1E2045", x"FFFDF6", x"FEFEFF", x"75719B", x"000F34", x"18334D", x"7797AE", x"000323", x"011C4E", x"071D41", x"041F47", x"0A1B47", x"000026", x"E3FCFA", x"FFF8EE", x"D4DDEB", x"051032", x"EFFDFF", x"FFF0FF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFF7F7", x"63728B", x"29345B", x"F6FFFB", x"FEFEF4", x"585E7C", x"050E39", x"031F3E", x"021C40", x"011C43", x"011C4A", x"2F3863", x"868B92", x"AEBFD9", x"00092F", x"0A1D42", x"0A1A54", x"A8AEC9", x"06092E", x"041F44", x"03214D", x"0C1F47", x"7684A3", x"FFFCF0", x"344270", x"FFF8FE", x"FDFFFB", x"FFFCFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFBF5", x"FAFFFB", x"5C6986", x"FBFEFA", x"3B5567", x"08214A", x"011B40", x"011B46", x"071E47", x"021B39", x"000020", x"A2A9BC", x"020E32", x"BBB9CD", x"DFF5E7", x"000B29", x"0C1C4A", x"0A2042", x"021D49", x"0A1D44", x"121C48", x"FFFFFF", x"FFFFF1", x"19294E", x"A4B1C4", x"FFF8FE", x"FFFFFA", x"F0FEF6", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"F9FFF5", x"FFFBFF", x"F8FBFF", x"121A3D", x"CACCDC", x"FEFCFF", x"CBCFD7", x"00042E", x"091B48", x"071E45", x"041F44", x"011B4A", x"7C8DA4", x"000021", x"022247", x"021D4E", x"000026", x"F5FFF9", x"3A5283", x"021C40", x"072046", x"011943", x"000031", x"F6FDFF", x"FEFFF1", x"01163D", x"FFFBFC", x"F9FEFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"F6FAFF", x"061746", x"FDFEEC", x"FAFFFF", x"02052C", x"071D4A", x"032048", x"0A1E47", x"071941", x"021D48", x"0A1F4D", x"000526", x"E8FFFF", x"101A49", x"09002E", x"02223B", x"021D42", x"021D46", x"021F43", x"383B60", x"FFFAFB", x"FAFFFC", x"01042E", x"FEFCFF", x"FBFEFA", x"F9FFF4", x"FCFBFF", x"FFFDF9", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFEFF", x"FAFFFB", x"FBFFF4", x"FFFEFA", x"97A8BC", x"3B4666", x"FFFFFC", x"F8FFF9", x"040020", x"0B214F", x"081F46", x"011C43", x"011239", x"011A4B", x"081C44", x"0B1940", x"A7C1D2", x"172B48", x"051A3C", x"011348", x"071F4C", x"021E3D", x"021D4B", x"11223B", x"FFFAFF", x"A8B6C9", x"E9F8F2", x"FFFEF9", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"E5F1FC", x"99AFBC", x"FDFEFF", x"0A1731", x"0A1F47", x"071D44", x"011C43", x"011942", x"051840", x"021B41", x"081C46", x"061C46", x"010E39", x"4E6385", x"0B1E47", x"011C43", x"081C44", x"041F45", x"3C4A63", x"FDFFF9", x"ECF2FA", x"1B264E", x"FFFEF5", x"FFFAFF", x"FCFCFC", x"FFFEFA", x"FFFCFF", x"FEFFFA", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FAFAFA", x"FFFFFA", x"FFFEFF", x"F5F6F0", x"F9FFF0", x"FEFEFF", x"020E32", x"FFFCFF", x"FAF6FF", x"020020", x"071948", x"021D41", x"072047", x"071F40", x"021B46", x"0B0A33", x"DFE5EC", x"000029", x"06133D", x"C3CED6", x"000326", x"021C42", x"061C46", x"05143C", x"DFE6F5", x"FFFAFA", x"011139", x"FFFEFB", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FEFFFF", x"FEFEFE", x"FEFDFA", x"FFF5F2", x"061638", x"FFF8FF", x"E8E4ED", x"01133D", x"021D42", x"061E4A", x"03143F", x"B4C0DB", x"96A5A8", x"34466D", x"051840", x"000233", x"324B78", x"041D42", x"061D44", x"021B44", x"0A1B50", x"242F4D", x"FFF3F5", x"D8F1E1", x"414B65", x"FCFBF9", x"FFFCFF", x"FAFFFB", x"FFFCFE", x"FFFBFF", x"FFFCFF", x"FFFCFE", x"FBFAF7", x"FBFFFC", x"FEF7FC", x"FFF2EA", x"FCFCFC", x"FFFFFC", x"FEFFFF", x"FFFFFF", x"F6FDFF", x"FFFFF4", x"F4F7FF", x"FFF8FF", x"FEFEFF", x"FFFFF6", x"F4FFFF", x"FFFCFF", x"FFFFFF", x"FFF4FF", x"FBFDF5", x"FEFEFB", x"FEFFFF", x"FEFFFF", x"FAFEFF", x"FFFAFC", x"FFFEFF", x"FFFEFF", x"F4FDFF", x"000527", x"FFFEFF", x"F6FFFE", x"00002C", x"062038", x"021F49", x"081B43", x"040C39", x"F1FEFF", x"668190", x"66748D", x"1F3557", x"07002C", x"1C4360", x"021E3F", x"022047", x"032439", x"0A0A36", x"FFFBFC", x"C2D1DC", x"E5EDF7", x"E9FFFB", x"FFFFFF", x"FFFDF9", x"FFFAF6", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFEFF", x"FEFDFA", x"F7F9FF", x"F3FFF5", x"8A9BA9", x"F4FFF6", x"081739", x"021F46", x"021C42", x"081F46", x"091C49", x"000C2A", x"374B72", x"8E9BB1", x"9C9FB5", x"FFFAF7", x"020825", x"0A1C45", x"021D4B", x"032145", x"000D32", x"F9FFFF", x"F4FFFF", x"2F416D", x"F8FFFA", x"FEFFF4", x"FFFEFF", x"FFFFFF", x"FFFFFF", x"061233", x"061233", x"061233", x"FFFFFF", x"061233", x"061233", x"F4FFFC", x"061233", x"F1F6F5", x"061233", x"EFF4F5", x"061233", x"F6FAFF", x"061233", x"ECF5EC", x"061233", x"061233", x"FEFEFF", x"ECEEE6", x"061233", x"061233", x"F7F8EE", x"061233", x"061233", x"F6FFFB", x"FFFEFA", x"F6FFF5", x"FCFCFF", x"FCFBF9", x"FBFFF1", x"F3FBFF", x"041133", x"FDFEF4", x"D4D8E4", x"0A0B40", x"011941", x"021F40", x"021E4C", x"011130", x"051B47", x"021C44", x"011A4E", x"011C47", x"0A2051", x"07133C", x"051B49", x"011C48", x"01163D", x"D3E5E8", x"FFFEFF", x"02164A", x"FFFBFF", x"FEFEF1", x"F5FFFF", x"FAFCFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFDF9", x"FFFBFC", x"F5FDF7", x"1B2B56", x"F3FFF4", x"FDEFF5", x"0A0E35", x"061D46", x"011941", x"011A3E", x"041E49", x"0D2050", x"375266", x"2E465E", x"022140", x"0E2C4D", x"021D4A", x"041D42", x"061E4A", x"000428", x"FEF9FA", x"F8FEF6", x"011132", x"FDFFF0", x"FFFFFC", x"FDFFFE", x"FEFFFF", x"FFFEF9", x"FEFFFF", x"061233", x"8297A4", x"F2FFF4", x"061233", x"F1FEFF", x"E0E8F5", x"061233", x"061233", x"F1FBFE", x"061233", x"F8FDFE", x"061233", x"061233", x"061233", x"FEFEFF", x"061233", x"FEFEFF", x"061233", x"FAFFFF", x"061233", x"F6FEFE", x"FDFFF1", x"061233", x"F1F9FF", x"061233", x"FBFCFF", x"FFF6F7", x"F7F7F7", x"FFFEFF", x"FFFFFC", x"FEFBFC", x"F8FFFF", x"3A4E6E", x"FFFCFF", x"5B7587", x"0C1A49", x"041F44", x"011B46", x"031B44", x"081B48", x"021D46", x"0A1439", x"000A2D", x"CDD0D6", x"818EA0", x"021F48", x"021D46", x"071E47", x"0C1948", x"F6FFF9", x"7890A1", x"FEFFFF", x"FCFAFE", x"F8FDFE", x"FFFEF7", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"F6FBFC", x"FEFFFA", x"F8FBFF", x"294064", x"FFFAFF", x"25395B", x"02224D", x"061B44", x"061D44", x"01143B", x"082148", x"071E49", x"011129", x"C2C3DF", x"132344", x"021D4A", x"081C44", x"092249", x"011640", x"AEBBDB", x"F2FFFF", x"000524", x"FFF3F7", x"FCF7FF", x"FFFFFF", x"FFFFFF", x"FEFEFB", x"FDFFFE", x"FBFFFF", x"061233", x"061233", x"E2E4E6", x"051A3C", x"FEFEFB", x"FFFCFE", x"061233", x"061233", x"FBFFFF", x"061233", x"FFFEFF", x"061233", x"061233", x"061233", x"FFFEFB", x"061233", x"FFFBFF", x"061233", x"FFFAFC", x"061233", x"061233", x"FFFDF6", x"061233", x"F9F5EF", x"061233", x"FFF7FF", x"FBF9FA", x"FFFFFF", x"F6F6F6", x"FEFEFF", x"FFFEFF", x"FFF9F1", x"AEB4C8", x"D5D9E7", x"FDFFF9", x"010B25", x"071A47", x"061D44", x"021D41", x"171E48", x"172F4D", x"DAD9E8", x"EEFDFA", x"0D172E", x"617790", x"00001C", x"031C45", x"011B40", x"090331", x"F9FCFF", x"FFFEEF", x"2F435F", x"FFFFFF", x"FFFDF9", x"FFFFF6", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FEFFFF", x"FAFFFC", x"96A9BA", x"FEFFF9", x"FFFBFF", x"000029", x"021C4C", x"0A1C47", x"06092A", x"6C7E98", x"090236", x"091F43", x"051D48", x"03223F", x"1B345A", x"031D40", x"021D4A", x"011C4D", x"031940", x"FFFEFF", x"7380A4", x"FAFFFF", x"FEFFFF", x"F1FAFF", x"FBFBFE", x"FAF8FF", x"FCFAFE", x"FFFCFF", x"FBFCFF", x"061233", x"60657E", x"FAFFFF", x"F4FDFF", x"061233", x"061233", x"F9FAFF", x"F6FBFF", x"061233", x"061233", x"FAFDF9", x"061233", x"F5FFFF", x"061233", x"F6FFFF", x"061233", x"061233", x"061233", x"EBF1EC", x"061233", x"061233", x"E4F9FF", x"061233", x"061233", x"F4FEFF", x"FBFFFF", x"FFFFFF", x"FFFEFF", x"FFFEFB", x"FFFEFF", x"FBFEF7", x"FFFFFA", x"FFFFFC", x"0A1739", x"FEFFF5", x"FEFFF5", x"090D2E", x"071845", x"0B1841", x"0A1541", x"E6EDFF", x"060A2D", x"000F34", x"4C5B7A", x"182145", x"415170", x"091C43", x"0C1C46", x"061A40", x"3A5879", x"FFFEFB", x"132B48", x"FFFAFF", x"FBFFFA", x"FDFEF6", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"F9FEFF", x"F8FDFE", x"0E254A", x"FBFCFF", x"A2B5CA", x"091B40", x"011A49", x"022045", x"17354E", x"CED0CD", x"FFFBFC", x"71848F", x"000F2D", x"415371", x"05133C", x"021F46", x"011C47", x"00082E", x"FFFBFF", x"F9FFF4", x"353F62", x"F9FDF1", x"FFFFF9", x"FFFEF9", x"FFFFFA", x"FFFFFA", x"FBFFFC", x"F9FEFC", x"FFFDF6", x"FBFFF6", x"FBFCFF", x"FFFFF4", x"F7F9F1", x"FEFFFF", x"FEFFFC", x"FEFFF5", x"FFFFFC", x"FEFFFA", x"F9FBF5", x"FFFFFC", x"FEFFF9", x"FFFFF9", x"FFFFFA", x"FEFFF7", x"F7F6F1", x"FDFFFE", x"FFFCFE", x"FFFAFA", x"FFFAF9", x"FFFBF9", x"FFFAEF", x"FFFFFA", x"FFFFFC", x"F6F8F0", x"FCFDFA", x"FFFEFF", x"FEFFFF", x"FEFFFC", x"FFFFFF", x"FFFFF9", x"FEFFFC", x"FFFEFF", x"FFFCFF", x"172D51", x"FFFAF5", x"284366", x"0A2048", x"022042", x"021E4A", x"021B38", x"1F354D", x"062D54", x"000B34", x"01183C", x"081C40", x"021B41", x"081B48", x"021D42", x"000028", x"F6FAEC", x"C3D4D7", x"E7E9F9", x"FFF6F2", x"F8FDFE", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFAF6", x"FFFEFA", x"364970", x"FFFCFF", x"13264A", x"022347", x"021D45", x"021F43", x"0A113D", x"0C1843", x"19354F", x"1A264A", x"F9FAFC", x"172E4A", x"021F4A", x"071E45", x"08214C", x"25375C", x"F5FFFA", x"132A51", x"F4FCEF", x"FEFAFF", x"FFFFFC", x"F5FCF6", x"FEFFFF", x"FFFBFC", x"FFFCFC", x"FFFEFF", x"FCFAFF", x"FFFFFC", x"FAFAFA", x"FFFCFE", x"FCFAFB", x"FFFBFB", x"FEF9FA", x"FFFFFF", x"FCFBF9", x"FFFCFF", x"FFFAFB", x"FAFAF7", x"FFFEF7", x"FEFBFF", x"FFFFF9", x"FFFCFF", x"FFFCFF", x"FFFFFC", x"FEFEFB", x"FFFFFF", x"FEFFFC", x"FEFEFF", x"FFFFFF", x"FEFFF9", x"FFFEFB", x"FFFFFA", x"FFFFFA", x"FFFFFA", x"FFFEFA", x"FFFEFC", x"FEFBFC", x"FEFEFF", x"FFF9FB", x"FAFFF7", x"FEFCFF", x"6E7F95", x"FBFAFF", x"FFF7FC", x"00012E", x"081C44", x"02234B", x"011740", x"5F7083", x"021739", x"011B48", x"071A46", x"000422", x"213762", x"011B45", x"041F44", x"0A0E3C", x"EAF0F5", x"FEFFFF", x"253E63", x"FFFFF9", x"F9FFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFAFF", x"B0C3CD", x"EBF1F6", x"FFFEFF", x"00002A", x"011A46", x"081E42", x"010C32", x"314A6E", x"0A0A39", x"7E9BB3", x"011948", x"021E3F", x"051A43", x"021C45", x"021C42", x"060E30", x"FDFEFF", x"F9FAFF", x"596C89", x"FEFEFF", x"FEFEFF", x"F7F9F1", x"FBFCFF", x"FBFDF5", x"FFFFFF", x"959EAB", x"9AABC7", x"9EAFBE", x"9DAFC3", x"9EAFC1", x"9CAEBF", x"97A8BA", x"A1B2C4", x"A0B1C3", x"A1AFC2", x"A0AFBE", x"A2B4C5", x"9AABBD", x"A3B2C2", x"A2B5C1", x"9FB0C2", x"9AADB8", x"9FB0C2", x"9EB1C2", x"9BADBE", x"9AABBD", x"A0B1C1", x"A3B1C4", x"9AA9B8", x"9FABC5", x"9DADBC", x"9FB0C4", x"97A8BC", x"9CAEC2", x"9BADBE", x"9CAFC4", x"98A2AE", x"FDFFF9", x"FFFFFA", x"FBFAFF", x"FCFAFB", x"FAFFF6", x"FFFBFE", x"0A2140", x"FFFEFF", x"213453", x"021E48", x"02203D", x"032146", x"203F6A", x"000020", x"192953", x"A4B7C3", x"FFF6FF", x"8F9BA1", x"081C44", x"021D45", x"041F47", x"465B83", x"FDFFFE", x"122C52", x"FFFFFC", x"FEFEFB", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFEF9", x"284168", x"FFFAFF", x"DDD9E5", x"021C40", x"021E4C", x"041F47", x"1A2E57", x"FDFFFB", x"FDF2F9", x"4B5D82", x"000129", x"1C2E5D", x"081A40", x"03244A", x"071A46", x"03153D", x"FEFEFB", x"243F67", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"596883", x"FFF8FE", x"EFF5F9", x"0B0D3C", x"032548", x"021E47", x"000025", x"FFF7FF", x"797E95", x"345070", x"000D38", x"617593", x"000929", x"021D42", x"011C42", x"040E38", x"F8FAF6", x"707C96", x"FFF9F6", x"FEFCFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FEF9F5", x"183157", x"FFFAFF", x"597088", x"071B45", x"041C43", x"031D40", x"0C2142", x"000F3B", x"000B2E", x"6D7189", x"FFF8FF", x"1A2944", x"0E1F53", x"051C42", x"081C44", x"98A7B1", x"FFFFF9", x"1F2F51", x"FFF7FF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"F6FFFF", x"425E7C", x"FBFFFF", x"000A33", x"021C3D", x"021C42", x"071A46", x"29415E", x"00113D", x"F6FFFF", x"93849B", x"FFFFFC", x"000B30", x"061F48", x"071A44", x"00012E", x"FEFFFA", x"F4FDFF", x"B5BFD4", x"FDFFFE", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFC", x"32476D", x"FCFBFF", x"0C2449", x"031C42", x"061C46", x"021F4A", x"0B1540", x"061D44", x"08143E", x"092541", x"213863", x"000C31", x"021E40", x"011B46", x"04082E", x"FAFCF4", x"D0CCE4", x"EAEEFC", x"FBFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FAFFF9", x"0E2552", x"FCFBF5", x"446580", x"062049", x"041F45", x"06204A", x"050030", x"FFF7FC", x"000024", x"00113B", x"00102A", x"071D47", x"021E46", x"091E48", x"06133D", x"DEE6ED", x"FFFFFA", x"2D476D", x"FDFFFB", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"F6FFFF", x"9EA4C1", x"FEFFFF", x"00032E", x"081B43", x"021A43", x"01133B", x"9D9EBC", x"1C3D5C", x"596587", x"100E36", x"01143F", x"011C49", x"071D41", x"051D48", x"0A1339", x"FFFBFF", x"183459", x"F5FCF6", x"FFFFFA", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFF5F9", x"8498AB", x"F8FFFF", x"DFE5EC", x"011439", x"061D46", x"051C43", x"05123B", x"304367", x"0A2246", x"081C46", x"031538", x"0C1A47", x"021D43", x"021E42", x"051A43", x"697D98", x"F1F1F4", x"193762", x"FFFCFE", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"ADB3CE", x"FBF6F5", x"FFFEFF", x"01012E", x"021F44", x"031D40", x"132240", x"152A4C", x"0B1646", x"7386A8", x"9197A9", x"6A7CA0", x"091B46", x"021F47", x"031C45", x"435A6C", x"FFFCFF", x"1D375B", x"FEFFFC", x"FFFFFF", x"FFFFFA", x"FCFBFF", x"FBFBF9", x"FFFFF9", x"FBFEF7", x"FCFDFA", x"FEFEFF", x"FFFCFE", x"FEFFF9", x"FFFFFF", x"FFFEFF", x"FFFCFF", x"FFFFF4", x"FFFCFE", x"FDFFFE", x"FEFFFF", x"FCF4FF", x"FFFDEE", x"FFFEFF", x"FEFEFF", x"FBFAF5", x"FEFCFF", x"FAFEF5", x"FEFFFF", x"F4FEFF", x"FCFBF5", x"FFF3FF", x"FFFBF7", x"FAFFFB", x"FAFEFF", x"FFF4F1", x"FEFEFE", x"FFFFFA", x"FEFFFF", x"FAFAFF", x"FFFAF6", x"F4FFF6", x"FAFBF5", x"FBFCFF", x"FFFFF6", x"FFFFF9", x"FBFFF1", x"FAFFFF", x"FFFFF9", x"FFF3FF", x"FFFFF6", x"798EAF", x"FEFBFC", x"02002A", x"021E43", x"021E3D", x"071B45", x"455880", x"3F4C6F", x"0B0331", x"FDFFF5", x"475570", x"0A1D4A", x"062141", x"021E4A", x"2B4B6F", x"FEF9F7", x"132E4E", x"FFFFFC", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"616F8F", x"FFFAFE", x"EBEFF5", x"02103B", x"0B1E51", x"021941", x"51657E", x"050034", x"0B1E47", x"011C52", x"00113B", x"7A91A1", x"021C46", x"021E48", x"071A44", x"A8B9C9", x"FFFFFA", x"4C6A7E", x"F9FBF5", x"FEFEFE", x"FEFEFF", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"F8FFFC", x"FBFEFA", x"061233", x"101E41", x"061233", x"061233", x"061233", x"FFFFFF", x"FFFAFF", x"F6FEFB", x"F1F6F7", x"FFFFFF", x"0F1940", x"082050", x"0D2142", x"000B39", x"FFFFFF", x"061233", x"061233", x"061233", x"061233", x"07163F", x"061233", x"F3FFFF", x"F3FBFF", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"FFFFFF", x"FEFAFF", x"F9FFF9", x"21375D", x"FAFAFC", x"031238", x"022047", x"061D40", x"000833", x"838CB5", x"011733", x"D8E2EB", x"001040", x"334F5B", x"02062D", x"031B49", x"091D41", x"0D2044", x"FCFCFF", x"3B587A", x"FDFEFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"385277", x"FFFBFF", x"B6C5CF", x"011845", x"072748", x"07214A", x"000B2F", x"6A798E", x"00012D", x"010C32", x"182448", x"2B4463", x"02224A", x"071E47", x"000F39", x"F6F7FC", x"DEE9E7", x"C0D5DA", x"FFFFF9", x"FFFFFF", x"FFFCFE", x"F9FEFC", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"FCF5F7", x"EDFDF1", x"061233", x"061233", x"061233", x"061233", x"FFFFFF", x"F6FFFF", x"FFF8FF", x"F9FDEF", x"061233", x"061233", x"061233", x"0B1A49", x"FFFFFF", x"FCFAFE", x"F9FFFF", x"061233", x"061233", x"061233", x"061233", x"FFFCFF", x"FFF9F9", x"FAF7FB", x"FFFFFA", x"061233", x"061233", x"061233", x"061233", x"FFFFFF", x"FFFFF1", x"FDFFFE", x"F3FFFB", x"183260", x"FFFFFF", x"1F375B", x"021C40", x"082043", x"0A1743", x"9BAFBD", x"3E4468", x"E9F8F7", x"00092B", x"BCD1EF", x"000E33", x"021E40", x"021E47", x"020B32", x"FFFEFF", x"6C809C", x"FAFBFE", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"16345A", x"FFFBFA", x"92A7AF", x"051947", x"071847", x"0A1E48", x"091D41", x"2C3750", x"FFFBFA", x"FCFAFF", x"A19DBD", x"07123C", x"011B48", x"021C42", x"000932", x"FFFEF7", x"8F9DB1", x"FBFFFF", x"FEFEF4", x"FFFFFC", x"FBFBFF", x"F9FFF7", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"FFF7F4", x"FEFFF9", x"061233", x"061233", x"061233", x"061233", x"FEFAFF", x"F1FDFB", x"F8FCFF", x"061233", x"061233", x"061233", x"12213E", x"FEFFF9", x"FFFEFC", x"FAFAFC", x"061233", x"061233", x"061233", x"061233", x"FFFCFF", x"FFFEFF", x"FBFFFF", x"FAF9F4", x"061233", x"061233", x"061233", x"061233", x"FFFFFF", x"FFFBFF", x"FFFFFF", x"FBFEFC", x"19345C", x"FFFFFC", x"4C6286", x"042046", x"021E42", x"021D45", x"0B0A40", x"0C2342", x"0B0838", x"041F48", x"01163C", x"0C1B4A", x"022141", x"031F4B", x"06002B", x"FEFAFF", x"A2A9BE", x"FFFEFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"183356", x"FAFBFE", x"798BA1", x"021F43", x"021A43", x"021C46", x"021D39", x"021E46", x"000428", x"00002B", x"0A1D48", x"031C47", x"021C46", x"031C42", x"000029", x"FEFBFC", x"5C7392", x"FEFEFE", x"FFFAF6", x"FBFEFA", x"FFFFFF", x"FDFFFE", x"000B39", x"061233", x"061233", x"000F31", x"FAFFFC", x"F9FFF9", x"FDFFFE", x"94A1B1", x"061233", x"061233", x"061233", x"061233", x"FEFCE9", x"FBFFFF", x"D5DDF1", x"061233", x"061233", x"061233", x"061233", x"061233", x"000929", x"061233", x"061233", x"061233", x"F3FFF5", x"FFFBFF", x"FFFBFF", x"FFFFFA", x"061233", x"061233", x"061233", x"061233", x"FBFFFF", x"FFFFFF", x"FFFCFE", x"FFFCFF", x"061233", x"061233", x"061233", x"061233", x"FFFFFF", x"FFFFFF", x"FFFEF7", x"FFFFFC", x"465A7A", x"FEFEFB", x"8190A8", x"031C47", x"021E46", x"051C43", x"162A52", x"000F3B", x"011139", x"011335", x"000A2B", x"172F4F", x"011B46", x"061E4D", x"00012B", x"FEFCFF", x"BDC8D0", x"EAEBF0", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"1A3659", x"FEFFFF", x"6E8096", x"022044", x"021F42", x"031B4A", x"374974", x"00052D", x"05002D", x"09002E", x"0B1536", x"08184D", x"021D47", x"071D44", x"00032D", x"FFFEFF", x"495F7C", x"FFFFFF", x"FFFDF9", x"FEFFFC", x"FFFFFF", x"FDFFFE", x"000B39", x"061233", x"061233", x"061233", x"FFFFF6", x"FFFFF0", x"FFFBFF", x"061233", x"061233", x"061233", x"00002C", x"FCFCFF", x"FBFFFF", x"FEFFF9", x"FEFDFA", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"F4FDF4", x"FFFEFC", x"FFFBFF", x"FFFFFA", x"061233", x"061233", x"061233", x"061233", x"FAFFFF", x"FFFFFF", x"FFFCFE", x"FFFCFF", x"061233", x"061233", x"061233", x"061233", x"FFFFFF", x"FFFFFF", x"FFFFF9", x"FFFFFC", x"556A8B", x"FEFEFB", x"8F9FB7", x"021B46", x"021E46", x"051C43", x"4E5B71", x"F4FFFE", x"FCFBFF", x"FFFBFF", x"FFFEFF", x"000E2A", x"0A1A4A", x"021C42", x"00012C", x"FEFCFF", x"CCD6DF", x"DADBE0", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"1B385B", x"FDFEFF", x"6B7D93", x"022045", x"021C41", x"0A1B43", x"909DAF", x"F9FEFF", x"FAFFF9", x"FFFCFF", x"F8FDFB", x"00021D", x"021E48", x"071D44", x"00032D", x"FFFCFE", x"475C79", x"FEFEFE", x"FEF9F5", x"FBFEFA", x"FFFFFF", x"FDFFFE", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"F9FBFF", x"F5FDF0", x"FAFFFF", x"FAFFF7", x"F8FDFB", x"FEFFFF", x"000025", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"FBF9FA", x"FCF6FF", x"FEFFFC", x"FFFBFF", x"FFFFFA", x"061233", x"061233", x"061233", x"061233", x"FAFFFF", x"FFFFFF", x"FFFCFE", x"FFFCFF", x"061233", x"061233", x"061233", x"061233", x"FFFFFF", x"FFFFFF", x"FFFFF9", x"FFFFFC", x"5B7193", x"FEFEFB", x"93A3BC", x"011B45", x"021D45", x"031C42", x"505E84", x"000020", x"070332", x"04012D", x"060022", x"2A3C6A", x"021D3F", x"021D43", x"02042E", x"FFFEFF", x"CFDAE2", x"D7D8DD", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"193558", x"FEFFFF", x"72849B", x"022044", x"092249", x"071D4B", x"283B63", x"000A33", x"02092E", x"050D33", x"001030", x"041F44", x"021D47", x"051C43", x"00012B", x"FFFEFF", x"526886", x"FFFFFF", x"FFFDF9", x"FEFFFC", x"FFFFFF", x"FDFFFE", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"FFFCFF", x"F4F6F5", x"FBFFFA", x"FBFAF7", x"FFFFF9", x"DFE7F4", x"061233", x"061233", x"061233", x"061233", x"061233", x"F9F9F9", x"FFFEF6", x"F8FFFC", x"F6FDF4", x"FFFBFF", x"FFFFFA", x"061233", x"061233", x"061233", x"061233", x"FBFFFF", x"FFFFFF", x"FFFCFE", x"FFFCFF", x"061233", x"061233", x"061233", x"061233", x"FFFFFF", x"FFFFFF", x"FFFEF7", x"FFFFFC", x"4C6182", x"FEFEFB", x"8797AF", x"031C47", x"021E46", x"051C43", x"011940", x"0A1F53", x"031E44", x"021E4D", x"0B1B41", x"061945", x"051C43", x"011B4D", x"00012B", x"FCFBFF", x"C4CFD7", x"E1E2E7", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"113457", x"FBFFFC", x"809BA0", x"071A49", x"081F46", x"082349", x"021B46", x"061C3E", x"011C43", x"091C4A", x"0E2940", x"0C2446", x"021F47", x"072047", x"00012E", x"FFFFF5", x"76859F", x"FAFAFF", x"FFFFF4", x"FFFFFA", x"FEFEFF", x"FBFEFC", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"FFFFFF", x"F6FFF6", x"F6FBFC", x"FFFEFA", x"FFFFFF", x"FFFFFA", x"061233", x"061233", x"061233", x"061233", x"061233", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FDFFF7", x"FFFBFF", x"061233", x"061233", x"061233", x"061233", x"FAFFFA", x"FCF8FF", x"FFFCFF", x"FFFFF4", x"061233", x"061233", x"061233", x"061233", x"FFFFFF", x"FFF6FF", x"FFFEFF", x"FFFEFF", x"2F4C73", x"FCFBF6", x"6F7CA4", x"022144", x"031E43", x"022046", x"01163B", x"081C4D", x"041C43", x"071643", x"828CAB", x"132A54", x"082045", x"071C43", x"090029", x"FEFAFF", x"ABB3C3", x"F5F5F5", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"1D3D60", x"FBFBFB", x"9AB4BB", x"011A47", x"021C42", x"011B43", x"081543", x"28365F", x"0A1942", x"00002A", x"FBFEFF", x"00012B", x"021F49", x"011B42", x"000B33", x"FFFEFC", x"B5C2C9", x"EAF5FB", x"FDFEF4", x"FFFFFF", x"FFFFFF", x"FDFFFE", x"061233", x"061233", x"061233", x"061233", x"FAFFF7", x"F9FFF1", x"FFF9F5", x"FAEFFF", x"061233", x"061233", x"061233", x"000A34", x"FEFFFF", x"FEF6F9", x"FFFBF7", x"FCFCFC", x"FFFEF9", x"061233", x"061233", x"061233", x"061233", x"061233", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFF7FF", x"FAFDF9", x"061233", x"061233", x"061233", x"061233", x"FCFBFF", x"FFFCEF", x"FAFBF5", x"FAFFFF", x"000C2A", x"061233", x"061233", x"061233", x"FFFFFF", x"FFFEFF", x"FCFCFC", x"FAFFFF", x"152F59", x"FBFBFB", x"304E6E", x"021F44", x"031D40", x"031B44", x"6E8CA9", x"00002F", x"00042A", x"040A25", x"465771", x"00082F", x"041D40", x"081B4B", x"02042E", x"FFFEFF", x"8696AE", x"FEFEFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"475F7E", x"FFFEFF", x"C6D5DC", x"011641", x"021C41", x"081E42", x"0A133B", x"ADB6C3", x"596D78", x"FBFFFF", x"04082E", x"071E49", x"021C46", x"021E46", x"01143B", x"DBE0EB", x"FBFFFA", x"8BA5B0", x"FDFFF9", x"FFFFFF", x"FFFFFF", x"FEFFFF", x"061233", x"061233", x"061233", x"091232", x"EBE7F5", x"F7ECF2", x"061233", x"061233", x"061233", x"061233", x"061233", x"0B1B3E", x"F8FFFF", x"FAFFFF", x"FFFAF6", x"FCFCFC", x"FFFFFA", x"061233", x"061233", x"061233", x"061233", x"061233", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFEFF", x"F4FEF0", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"FDFFFE", x"FFFCFE", x"FEFEFF", x"F0FEF6", x"1D3561", x"FFFFFF", x"0D2646", x"031E46", x"081E42", x"01143E", x"C5DBE2", x"FFFCFF", x"FFFEF5", x"FBF6F2", x"F0FAFE", x"05002F", x"0A1F4A", x"021B44", x"061439", x"FBFCFF", x"587192", x"FEFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"838FAB", x"FEFEFE", x"F9FEFF", x"010A32", x"061D4A", x"03203D", x"2C3D71", x"00002A", x"060027", x"5E6983", x"56628C", x"718BA5", x"031D48", x"021D46", x"061B44", x"708795", x"FCFAFB", x"26415F", x"FAFDF6", x"FEFEFE", x"FEFEFF", x"F9FBFA", x"061233", x"061233", x"061233", x"061233", x"041039", x"09103D", x"061233", x"061233", x"061233", x"061233", x"061233", x"FFFFFF", x"FAFFFA", x"F6FFFF", x"FFFDF9", x"FEFEFE", x"FFFEF9", x"061233", x"061233", x"061233", x"061233", x"061233", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"F9FBF7", x"F9FEFC", x"FCFAFB", x"040323", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"040024", x"FFF8FF", x"F7F6FE", x"FCFDFA", x"FFF8FF", x"FBFFF4", x"3B5070", x"FFFEFF", x"00052F", x"022248", x"041E3F", x"051A43", x"011938", x"01143D", x"001034", x"00012E", x"787E8B", x"001139", x"0B2045", x"051D48", x"1B3357", x"FFFEFF", x"234064", x"F4FBF9", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"D3E2DC", x"DAD9E8", x"FBFFF4", x"04002A", x"022045", x"021F44", x"00001D", x"FAFFFF", x"E7E8EB", x"727E9B", x"2C3367", x"7D95A9", x"051940", x"061F48", x"081C43", x"213961", x"FFF7F7", x"0F2C56", x"FDFEFF", x"F9FFF9", x"FFFFFF", x"061233", x"00001C", x"04012D", x"02002D", x"02002D", x"02002D", x"02002D", x"061233", x"061233", x"061233", x"182A45", x"FFFFFF", x"FBFEFC", x"FFFFFC", x"FFFFFF", x"FBFBFB", x"FBFEF7", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"FAFDF9", x"FFFFFA", x"FFFEFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"061233", x"F7F6FC", x"FAFAFC", x"FEFEFE", x"FFFFFC", x"FFF7F9", x"D9DADF", x"DAE6F2", x"F8FFFF", x"00032F", x"022141", x"022049", x"051D48", x"021B44", x"021D40", x"031F41", x"021137", x"F2FFFF", x"051446", x"071A47", x"021D4A", x"4B5D7F", x"F8FFFF", x"1B2E5C", x"FCFCFC", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"F9FFFA", x"667693", x"FCFCFC", x"011039", x"021E43", x"011C43", x"04123D", x"192B4D", x"0A1940", x"021F43", x"000D34", x"070738", x"071D43", x"071E49", x"051B45", x"00012D", x"FFFBF9", x"5D7493", x"FAFFFF", x"FBFAF5", x"FFF8FE", x"F7F9FE", x"FEFEFF", x"FFFEFF", x"FEFCFF", x"FEFCFF", x"FEFCFF", x"FEFCFF", x"F6FEFE", x"FAFFFF", x"FFFFFF", x"FFFEF7", x"FFFFFF", x"FFFFFC", x"FFFFFC", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FBFFFF", x"F6FFFF", x"FCFAFB", x"FFFFFC", x"FBFEF7", x"FAFDF6", x"FBFFFF", x"F9FBF7", x"FEFEFB", x"FCFCFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FAFFFB", x"F9FEFF", x"FEFFFF", x"FAFBFE", x"FAFAFA", x"FFFFFF", x"FFFFFC", x"FBFFF4", x"FBFBFE", x"FFFFFF", x"FFFFFF", x"FFFFFC", x"FEFFFF", x"284569", x"FBFAF5", x"9FB0C2", x"071B45", x"0A2048", x"011C48", x"01193A", x"031E43", x"032146", x"022047", x"022249", x"000A29", x"02224B", x"031D40", x"021742", x"A3B5C7", x"FFFFFA", x"213865", x"FCFDFA", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFEFC", x"223C61", x"FFFCFF", x"244162", x"021C44", x"041F45", x"021D42", x"071E47", x"0A1548", x"0A082F", x"FBFEFC", x"F0EDF4", x"000625", x"0B1E4A", x"021F48", x"021039", x"EFFAF4", x"FFFBFF", x"75819C", x"FBFCFF", x"F7F9FB", x"FEFFFF", x"FEFEFB", x"FEFDF7", x"FFFEFF", x"FFFEFF", x"FFFEFF", x"FFFEFF", x"FAFAF7", x"FFFFFF", x"FCFCFC", x"FFFFFF", x"FCFDFA", x"FFFFFA", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFCFE", x"FEFDFA", x"FEF7FC", x"FFFAFF", x"FFFCFF", x"FFFFFF", x"FFFFFF", x"FBFBF9", x"FFFFFF", x"FCFCFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFCFC", x"FEFDFA", x"FAFFFF", x"F5FAFF", x"F4FFFF", x"FAFFFF", x"FBFCFF", x"FFFFFF", x"FFFFFF", x"FCFCFC", x"FEFEFE", x"FFFFFF", x"F5FEF5", x"132855", x"FEFEFE", x"122C4F", x"091C49", x"021B41", x"06224B", x"3F4F6E", x"000B31", x"0A1D46", x"040F33", x"040926", x"34486C", x"06204A", x"0A1947", x"000D34", x"F4FFFB", x"FCFCFC", x"5D7191", x"FFFFFC", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFEFF", x"12284F", x"FFF6FF", x"9AA1B6", x"081F46", x"011B42", x"082043", x"0A1440", x"BFD4D4", x"A7B2BE", x"1A365B", x"00021C", x"6F7EA5", x"0A1D46", x"021D47", x"011B40", x"3D4F6F", x"F6FDF4", x"061B3B", x"FFF8FF", x"FAFFFF", x"F3FAFA", x"F9FFFF", x"F8FFFF", x"FFFFFC", x"FFFFFC", x"FFFFFC", x"FFFFFC", x"FAFFFB", x"FEFFFC", x"FEFEFB", x"FFFEFF", x"FEFBFC", x"FEFBFC", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FEFEFE", x"FFFCFF", x"FEFEFF", x"FAFAFC", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FAFAFA", x"FEFEFE", x"FFFFFC", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FBFEFA", x"FEFFFC", x"FCFDFA", x"FDFEF7", x"FFFEFF", x"FEFEFF", x"FBFBFB", x"FEFFFF", x"FCFDFA", x"FBFBFB", x"FFFFFF", x"FBFBFB", x"DEECFE", x"CBDBE8", x"F5FBFF", x"00002F", x"022047", x"021D40", x"000931", x"F0FBFF", x"FBF9FC", x"83808C", x"FBFBFF", x"FEFFFF", x"000029", x"021F41", x"032045", x"000029", x"FEFFFA", x"B2BED5", x"F1EEF5", x"FBFAFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FCFAFE", x"5E7F88", x"FFFCFF", x"F6FAFF", x"0B0A32", x"071F4E", x"021E3E", x"00002A", x"687891", x"000613", x"2F4765", x"A6AECA", x"F9FCFF", x"01112E", x"011A44", x"021C42", x"000226", x"FFF5F9", x"BBB5C7", x"F0FAFE", x"FEFFF2", x"FDFFF9", x"FFFFFF", x"FEFFFC", x"FCFCFC", x"FBFFFF", x"FEFFFC", x"FFFFF9", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"F9F9F6", x"FEFBFC", x"FEFBFF", x"FEFBFF", x"F9FFF1", x"FFF9F9", x"F1F9EC", x"FFF8FF", x"091C3D", x"F6F3FA", x"8B9EAC", x"031D48", x"041F48", x"062049", x"0B214B", x"00113A", x"02002A", x"8C9BC2", x"000015", x"011142", x"0A1C48", x"021C3C", x"021843", x"1B3062", x"FBFEF7", x"2D4867", x"FFFEFB", x"FFFCFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFF6FF", x"F9FEFF", x"A2AFBD", x"FDFEF7", x"000A2E", x"04214A", x"051C42", x"01153B", x"C8D1E1", x"FFF4FF", x"AEAEBA", x"071941", x"071033", x"0A1D48", x"021B44", x"092046", x"031F41", x"97A9BD", x"F2FFFE", x"011740", x"FBFFFC", x"FFFCFF", x"FFFFF6", x"FEFFFF", x"FBFBFB", x"FCFBF5", x"F8FAF6", x"F4FFFE", x"FEFFFF", x"FEFFFF", x"FEFFFF", x"FEFFFF", x"FEFFFF", x"FEFFFF", x"FEFFFF", x"FEFFFF", x"FEFFFF", x"FEFFFF", x"FEFFFF", x"FEFFFF", x"FEFFFF", x"FEFFFF", x"FEFFFF", x"FEFFFF", x"FEFFFF", x"FEFFFF", x"FEFFFF", x"FEFFFF", x"FEFFFF", x"FEFFFF", x"FEFFFF", x"FEFFFF", x"FEFFFF", x"FEFFFF", x"FEFFFF", x"FEFFFF", x"FBFBF9", x"FFFEFB", x"FFFEFC", x"FFFCFB", x"FFFBFF", x"FBFFFC", x"F5FDF7", x"FFFFFF", x"7F8BB0", x"F6FEF9", x"060434", x"011A47", x"061D46", x"031E46", x"031C45", x"0A1E49", x"071F42", x"000B2F", x"BDC0D5", x"233D5F", x"021F44", x"081E45", x"061C4A", x"93A3BA", x"FEFFFF", x"112A56", x"FEFFFA", x"F8FDFB", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FBFBF9", x"FCFAFE", x"162E58", x"FFFFFC", x"455B7B", x"041D42", x"031C47", x"022247", x"4F6591", x"000226", x"021C42", x"011843", x"081E4A", x"021D41", x"021C42", x"051B45", x"051A4A", x"00002D", x"FFF9F9", x"AFC0D2", x"E1ECF2", x"FFFCFE", x"FCFBF9", x"FEFFF7", x"FFFFFC", x"FEFFFF", x"435065", x"465F86", x"485F7E", x"485F7E", x"485F7E", x"485F7E", x"485F7E", x"485F7E", x"485F7E", x"485F7E", x"485F7E", x"485F7E", x"485F7E", x"485F7E", x"485F7E", x"485F7E", x"485F7E", x"485F7E", x"485F7E", x"485F7E", x"485F7E", x"485F7E", x"485F7E", x"485F7E", x"485F7E", x"485F7E", x"485F7E", x"485F7E", x"485F7E", x"485F7E", x"4A6086", x"424F66", x"FAFFFF", x"FFFEFF", x"FFFFF9", x"FEFFF9", x"FFF6FE", x"011537", x"FFFFFC", x"B3C3D2", x"031D40", x"021E42", x"011A42", x"071E47", x"021C44", x"021C44", x"061945", x"0B1D49", x"323D5F", x"050E3A", x"091A47", x"021D47", x"00002E", x"FFFFF4", x"F8FEF6", x"70809D", x"FFFEFA", x"FAFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FAFFFE", x"F8FCFF", x"253D5B", x"FFFEFB", x"EBF0FB", x"051034", x"031D4D", x"011B43", x"031439", x"022047", x"011B45", x"032545", x"091F47", x"041F45", x"0A234B", x"041F45", x"021E48", x"041F45", x"869BB4", x"FFFEF2", x"05092D", x"FBFFFA", x"FCFBF6", x"FEFFFF", x"FEFFFF", x"FCFAFE", x"FFF8FF", x"FFF7FF", x"FEFFFC", x"FEFFFC", x"FEFFFC", x"FEFFFC", x"FEFFFC", x"FEFFFC", x"FEFFFC", x"FEFFFC", x"FEFFFC", x"FEFFFC", x"FEFFFC", x"FEFFFC", x"FEFFFC", x"FEFFFC", x"FEFFFC", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FEFFFC", x"FEFFFC", x"FEFFFC", x"FEFFFC", x"FEFFFC", x"FFFFFF", x"FEFFFF", x"F9FFFA", x"F9FFFB", x"F8FAF9", x"FCFAFB", x"BFCBE2", x"C0D5E6", x"FBFFF9", x"000027", x"011B46", x"061B41", x"062049", x"011B43", x"031C45", x"021D45", x"031D40", x"011D51", x"01183E", x"072049", x"051D48", x"021A43", x"141D3E", x"FEFFFC", x"617A90", x"FFFBFF", x"F9F8F2", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"F8FEFF", x"FBFFFC", x"F5F3FF", x"A2C5CE", x"FBFCFF", x"020F30", x"031844", x"031F41", x"021D45", x"021E46", x"021C44", x"061D46", x"021E40", x"0A1844", x"071F44", x"021E40", x"031E44", x"022047", x"000928", x"FFFCFF", x"F4FFFE", x"38526A", x"FEFFFC", x"F9FFFF", x"FDFFFB", x"FFFEFB", x"FFFFFC", x"FAFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FEFEFE", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FBFEF7", x"FBFEFC", x"FFFFFC", x"FEFEFB", x"FFFAFF", x"051939", x"FFF3F7", x"6C798E", x"0A2149", x"031C41", x"011B45", x"021C46", x"051947", x"022247", x"011B46", x"071D47", x"031C45", x"021B44", x"022047", x"02204B", x"021D45", x"9FB8CE", x"FFFBF7", x"0D2147", x"F9FAF2", x"FFF9F5", x"FAF8FF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FEFDFA", x"FBFFFC", x"0B1A4A", x"F9FBFA", x"8993B0", x"071D44", x"031F47", x"031E46", x"021D45", x"031E46", x"071E47", x"071739", x"00082E", x"091F49", x"03204A", x"041C43", x"051B45", x"051A4A", x"1B224A", x"F9F9FF", x"9C9CB6", x"D4DFE5", x"FFFAFC", x"FBF8FF", x"FEFCFF", x"FFFFFF", x"FFFFFC", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"F9FFF5", x"FFFFFF", x"FAFFFF", x"FFFFFF", x"061233", x"FCFBFF", x"F9FFFA", x"FFF6EE", x"FFFCFF", x"FFFEF7", x"FFFCFF", x"FBFAFF", x"FFFFFF", x"FEFEFE", x"FFFFFF", x"FCFCFC", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFC", x"FFFFFF", x"FFFCFF", x"FFFEFF", x"FAFFF5", x"00072B", x"FDFDF2", x"F0FFF7", x"00012B", x"021A4A", x"021E41", x"021C46", x"0A1D43", x"011746", x"01002E", x"061E4B", x"021D45", x"021E46", x"081B45", x"021A43", x"0C1F48", x"000029", x"FFFEF5", x"FEFFFC", x"9CA8BF", x"FBFBF9", x"FEFFFF", x"FEFFF6", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFBFC", x"FFFFF9", x"F6FBFC", x"748A9F", x"FFFFFF", x"FFFEF0", x"000029", x"081C46", x"021D45", x"021E46", x"061D46", x"011740", x"E6E3F5", x"FFF3F9", x"000026", x"032348", x"021B44", x"022043", x"061C46", x"0D1A45", x"8BABB4", x"FFF7FF", x"1B3557", x"FFFBFF", x"FDFEF6", x"FEFFF9", x"FEFCFF", x"FEFDFA", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"061233", x"FFFFFF", x"F4FFF5", x"19284D", x"FFFFFF", x"061233", x"FFFFFF", x"061233", x"061233", x"FBFFFF", x"061233", x"061233", x"FAFAFA", x"FEFEFE", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFEFF", x"FEFEF1", x"FDFFFB", x"2C3963", x"F4FFFF", x"FFFAFF", x"000129", x"061D44", x"042247", x"051A40", x"061D4A", x"08194B", x"50608D", x"FFFEFB", x"011739", x"081B45", x"021D45", x"021B44", x"021F46", x"022249", x"4F678A", x"F1F9F9", x"122B55", x"FFFCFB", x"FFFFFC", x"F8FEFF", x"FEFEFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFC", x"FCFCFC", x"FFFEFF", x"FFFFF1", x"203652", x"FBF9FC", x"557086", x"061E4B", x"021C44", x"041F47", x"061C46", x"01163E", x"6F7896", x"D2D1F5", x"020F38", x"022047", x"031E46", x"071B45", x"022245", x"041F45", x"000430", x"EDFAF2", x"FFFCFC", x"01112E", x"F5FFFF", x"FDFEF6", x"FAF7FE", x"FBFEFA", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"061233", x"FFFFFF", x"FFFFF6", x"FFFFFF", x"061233", x"FBFFFF", x"FFFFFF", x"F3FFFF", x"061233", x"F3FFF9", x"061233", x"FFFCFE", x"FFFFFF", x"FEFEFE", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"F7F6F4", x"F5FDF7", x"616A87", x"E0E3EC", x"EDF9FA", x"16244E", x"021C42", x"051C42", x"031E44", x"041F47", x"021F44", x"021B44", x"0D1E40", x"E9F4FA", x"30416A", x"081B45", x"021C44", x"031C45", x"021D45", x"000029", x"FAFFFA", x"FFFBFF", x"3F4A6E", x"F3FFF5", x"FFFFFF", x"FDFFFE", x"FFFEFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"3F5B84", x"FFFFFC", x"FDFEFF", x"000226", x"091B43", x"031E43", x"051B47", x"011B45", x"031C45", x"01153D", x"091F49", x"031E46", x"011A40", x"071A4A", x"031A3E", x"081B4A", x"021E46", x"000028", x"FFF4FF", x"F3FFEB", x"090F2F", x"EEFFFF", x"FFF8FF", x"F6FFFF", x"FFFEFF", x"FEFFFA", x"FEFFFA", x"FFFFFA", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"061233", x"FFFFFF", x"FFFFFF", x"061233", x"F6FFFF", x"061233", x"FFFFFF", x"061233", x"F3FEFA", x"FFFAFC", x"FFFFFF", x"061233", x"FFFFFF", x"FEFEFE", x"FEFEFE", x"FFFFFF", x"F9F9F9", x"F9FAFC", x"FEFFFA", x"FFFBFF", x"FDF3FF", x"F9FBF7", x"494F74", x"D6DAE5", x"FFFFFC", x"4E5577", x"081C44", x"011C43", x"02174D", x"031940", x"021E40", x"021B44", x"021B44", x"061B44", x"01133A", x"051B45", x"041F4A", x"071A42", x"0A2447", x"031F47", x"435978", x"F8FFF2", x"313F62", x"FFFDF6", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFC", x"183157", x"FFFEFC", x"74879F", x"022044", x"022145", x"031E46", x"031E46", x"011B42", x"071E47", x"021C44", x"031F47", x"061847", x"112545", x"011A47", x"022049", x"061D46", x"091B43", x"000721", x"FFF7FF", x"FEFFFF", x"272A59", x"CDD9D7", x"F5FAFB", x"FAFBF5", x"FFFFFF", x"FDFEF4", x"FEFBFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"061233", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"061233", x"F3FEFA", x"FFFFFF", x"061233", x"FFFFFF", x"FEFFFF", x"FAFFFF", x"061233", x"FFFFFF", x"FEFEFE", x"FEFEFE", x"FEFEFE", x"FFFFF9", x"FBFBFB", x"FFFFF9", x"FFFEFF", x"F5FFF4", x"141E44", x"EFFAFF", x"FFF5FA", x"5C687C", x"021B37", x"011B43", x"081B43", x"021B3F", x"011439", x"022049", x"021E3F", x"021C44", x"061D46", x"071E47", x"021D45", x"021E44", x"022047", x"071641", x"00042B", x"FFFBFE", x"FFFDF9", x"364D68", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FDFEFF", x"66768F", x"FAFFF6", x"FFFFF9", x"050022", x"021843", x"08214A", x"011942", x"041F48", x"021C44", x"041F47", x"011B43", x"0A214A", x"0F1038", x"5E7985", x"071940", x"021B44", x"021D47", x"0A1D46", x"000028", x"EEF0EC", x"F9FAFF", x"8C91AD", x"454B67", x"FAFFFF", x"FEFEFB", x"FFFBFF", x"FAFEF5", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FAFBFF", x"FFFFFF", x"FFFFFF", x"FEFFFC", x"FBFFFF", x"FCFBFF", x"FFFFFF", x"FEFFF5", x"FFFFFF", x"FFFFFF", x"061233", x"FEFBFC", x"FEFEFE", x"FEFEFE", x"FFFFFF", x"FFFFFF", x"FBFCFF", x"FFFBFF", x"FAFEF5", x"F4FEFF", x"010826", x"F9FFF9", x"FFFCFF", x"314060", x"071D41", x"071E47", x"0A1A48", x"021C40", x"000A32", x"7F89A9", x"011746", x"022044", x"021E46", x"021C44", x"031E46", x"021E46", x"021C42", x"051D48", x"0C2149", x"8FA0BE", x"F6F5FC", x"172E58", x"FFFFF9", x"FBF9FC", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFF9F1", x"FFFFFF", x"000C34", x"F9FEFC", x"DCE6F6", x"000E36", x"051C43", x"021E4A", x"031E46", x"031F47", x"031C45", x"071B45", x"00092B", x"FFFAFF", x"1B1F34", x"303D60", x"011940", x"031C45", x"021B44", x"031F47", x"000B35", x"8599A4", x"FDF2FF", x"F6FFFF", x"060A29", x"E9EAFA", x"FEFFF9", x"F8FEF6", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FEFDFA", x"FBFDF5", x"FFFFFF", x"FFFEFF", x"F9FDEF", x"FEFFFF", x"FEFFF9", x"FFFCFB", x"FEFEFE", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFA", x"F6FAF1", x"4B4D71", x"556386", x"FAFEFF", x"FEF7F2", x"02103B", x"021A45", x"081B45", x"021C44", x"0A1C45", x"09163E", x"6B729A", x"FCFAFB", x"000A29", x"0B1E47", x"021D45", x"061D46", x"021B44", x"021D45", x"091A45", x"071941", x"0A0E2A", x"FFFFFA", x"F3FFFF", x"8291A7", x"FAFEF2", x"FBFBFB", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FCFCFC", x"FDFFFB", x"E7E4F5", x"98B2D4", x"F9FFF5", x"3A4866", x"08214C", x"022349", x"031B44", x"051746", x"11244B", x"0F143A", x"FEFAFF", x"020525", x"00011F", x"F6FFFB", x"011937", x"09203F", x"011B51", x"03244A", x"011B41", x"021B44", x"1F274A", x"FFF4FF", x"FDFEF4", x"9FABBC", x"111A44", x"EAF6F7", x"FEFFFF", x"FFFEFF", x"FCFDFA", x"FEFFFF", x"F4F9F7", x"FDFFFE", x"FFFFFC", x"FFFFFF", x"FDFFF9", x"FEFFFA", x"FEFFFA", x"FDFFF9", x"FDFEF7", x"FDFFFE", x"FEFFFF", x"F9FEFC", x"FEFFFF", x"FFFEFB", x"FBFBFE", x"FBFEFC", x"6D7893", x"17234A", x"F8FFF6", x"FFF7FF", x"B8BAD6", x"000628", x"071F44", x"021F46", x"02234B", x"0A1E46", x"01093F", x"26435E", x"03153D", x"00021B", x"F8FEF6", x"07052F", x"0A1947", x"022040", x"08184A", x"011B45", x"091F46", x"00002B", x"FBFFFF", x"FFFDF7", x"000324", x"FFFFF9", x"F4F9FC", x"FFFBF7", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FCFDFA", x"FAFDFB", x"FDFEF7", x"222E4B", x"FEF7F4", x"F8FCFF", x"000021", x"0A1E3F", x"071C42", x"071D44", x"071A30", x"FFFEF9", x"00012A", x"344F6C", x"EBEAFA", x"04102B", x"0C1741", x"394E6E", x"011240", x"021D3D", x"011940", x"021843", x"0A214C", x"000527", x"8995AE", x"FFF6F5", x"F8FFF9", x"A2A7BD", x"12183F", x"868D9F", x"FEFFF6", x"FEFFFF", x"FBFFFF", x"F9FFFA", x"F9FDF4", x"FAFEF2", x"FFFFFA", x"FEFFF9", x"FFFFFA", x"FFFFFA", x"FBFFF4", x"FDFFF9", x"F9FEFC", x"FAFFFE", x"F8FAF4", x"E6EEEB", x"313757", x"232D59", x"F9FCFF", x"F9FFF6", x"FFFBFF", x"1B2245", x"011139", x"061A48", x"081F48", x"011944", x"091C43", x"00113A", x"C5E5F0", x"5A6A7C", x"00052A", x"B1CCD5", x"00041C", x"FFFEFC", x"939BB4", x"000F36", x"03234A", x"022044", x"071D49", x"869AA7", x"FEFFFF", x"535D7E", x"F4FFFF", x"FFFCFF", x"F6FBFA", x"FEFDF6", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FCFCFF", x"FFFFF9", x"FEFEFF", x"F6FFFF", x"000527", x"FBFFFF", x"F6FDFF", x"000126", x"071843", x"011B42", x"0A1E4F", x"13294E", x"01173C", x"061A46", x"011642", x"041E4D", x"000027", x"FAFDFB", x"8B9FAF", x"000B3C", x"021D43", x"051C43", x"022042", x"0A1A46", x"082043", x"02002C", x"96A2B3", x"FFFBFF", x"FEFEFB", x"FEFFFF", x"566082", x"111E4A", x"314362", x"9BABB5", x"F2F4F6", x"FFFBFF", x"FAFFFF", x"FAFFFF", x"FAFFFF", x"FAFFFF", x"FFFCFF", x"CCD5D9", x"6C7E94", x"203155", x"1D2A51", x"ABB1C4", x"FFFFFA", x"FCFDFA", x"FBFAFF", x"364367", x"00002B", x"09234B", x"0A2048", x"021D40", x"021C40", x"011B41", x"011842", x"0C214A", x"00022A", x"BECED9", x"C8CEE2", x"040028", x"031D4A", x"5C7691", x"000025", x"081E4A", x"022042", x"061E4A", x"173049", x"FCF7F6", x"FBFBFF", x"717E93", x"FFFEFF", x"FBF6F7", x"FCFDFA", x"FBFDF5", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FBFDF6", x"FFFEFF", x"FFFFFA", x"FEFEFB", x"FAFFFF", x"475972", x"FCFCFC", x"B8D1DF", x"011134", x"061B44", x"02203F", x"021D47", x"0A1942", x"061C40", x"062045", x"000126", x"FDFFF7", x"060320", x"04022B", x"6B859D", x"021B44", x"061D46", x"021E40", x"031E46", x"021D45", x"061D4A", x"031C3D", x"00002C", x"455372", x"EBEEEC", x"FFFAFA", x"FFFFFA", x"FAFDF9", x"F4FFF5", x"AFC0C3", x"66778C", x"49607D", x"3C516E", x"415774", x"4F6684", x"7E8F9D", x"D5E4DF", x"FBFFFA", x"FEFEFF", x"F7F6F4", x"FEF9F5", x"ABB6C1", x"0A173A", x"000B2F", x"021F47", x"011845", x"071D49", x"061E4A", x"011C43", x"031843", x"011130", x"022047", x"022044", x"061B44", x"000737", x"AFCCD0", x"666A90", x"243860", x"031342", x"021F44", x"021D45", x"051B47", x"02002C", x"FBFCFF", x"FFFAFA", x"060F36", x"FCFCFC", x"FFFFFF", x"FEFFF6", x"FFFFFA", x"FFFEFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FDFEF4", x"ABAECF", x"C4C7DA", x"FFFFF0", x"7C8E9E", x"061A3C", x"031B44", x"021E4A", x"022045", x"011941", x"0A2046", x"DBE6FB", x"2D344D", x"7C93AB", x"FFFCFF", x"18214C", x"042042", x"022248", x"031647", x"041D4C", x"091A49", x"022349", x"07174A", x"021F40", x"091F46", x"090E39", x"00012E", x"1D3755", x"8490A3", x"DCE6F2", x"FEFFFF", x"FFFFF9", x"FFFEFF", x"FFFCFE", x"FFFEFF", x"FFFCFE", x"FEF9FA", x"FAFBFF", x"BAC8D6", x"576977", x"091235", x"00002B", x"081C46", x"041C43", x"021B44", x"03204A", x"082045", x"0A174C", x"011A3A", x"022045", x"011339", x"FFFEF9", x"404A64", x"011039", x"091B46", x"021D42", x"00002A", x"FAF4FF", x"01002D", x"011C43", x"021D4D", x"0B1E3E", x"000027", x"F4FFF7", x"FFFEFF", x"00041C", x"F9FFF6", x"FFFEFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFF6", x"FCFBFF", x"455672", x"E9FFFF", x"FFFEFC", x"567585", x"051A43", x"051745", x"021B44", x"0A1E4A", x"171C3D", x"EFEEEB", x"0E0027", x"FDFDEE", x"000028", x"041F45", x"050D33", x"627198", x"72829C", x"657994", x"01012F", x"071C43", x"011B3C", x"022046", x"021D41", x"022144", x"061D4A", x"021B46", x"061B42", x"06133B", x"02052C", x"090029", x"00012C", x"050830", x"02052E", x"00002A", x"000026", x"060D34", x"06153E", x"0A1E49", x"071D49", x"022044", x"042046", x"021D41", x"021E48", x"081F46", x"0A1E4A", x"000326", x"91A9C2", x"00002C", x"061943", x"58768B", x"4D5A78", x"F1EFF2", x"00002C", x"000F3F", x"0B244A", x"06173A", x"031C47", x"021E40", x"031C45", x"00012A", x"FEFAFF", x"FFFEF2", x"101D46", x"F6FFFF", x"FBFAF5", x"FEFCFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFF0", x"FFFFFF", x"1D254E", x"F5F9FF", x"FFF6F9", x"507384", x"02143B", x"011B40", x"022042", x"021C44", x"04123D", x"010529", x"E2DBF5", x"031E4A", x"09163E", x"D0DFDC", x"121E3C", x"021B39", x"000020", x"FFFAFF", x"021241", x"011443", x"021F3E", x"071A46", x"021C43", x"082147", x"031C45", x"091A45", x"011C47", x"011B4A", x"0A1C4D", x"051C43", x"051C43", x"051C43", x"031C42", x"0A1D4B", x"011C48", x"071E49", x"091A47", x"071F44", x"041F44", x"021D43", x"071845", x"01193D", x"000028", x"7D89A1", x"8E92AC", x"00092D", x"11284E", x"051743", x"506377", x"688197", x"0B0D34", x"F6FFF9", x"6D7893", x"01113F", x"022045", x"061F48", x"071E47", x"000024", x"FFFBFF", x"FEFFF6", x"273966", x"F8FEF9", x"FFFFFA", x"FFFEFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FDFEFF", x"FBF9FC", x"F9F6FC", x"FBFFEA", x"111B45", x"F6FAFF", x"FEFDF7", x"738494", x"020D37", x"051D48", x"051842", x"021E42", x"091B46", x"98A6B0", x"011235", x"0A0029", x"FFFFF9", x"040139", x"011A42", x"011B49", x"9AABB0", x"031332", x"203B5A", x"6E7D96", x"203759", x"021A43", x"01153A", x"051A43", x"021F46", x"061B44", x"061C46", x"021D44", x"021E48", x"021E48", x"021E48", x"021C46", x"021C44", x"061D46", x"021D45", x"022147", x"011C43", x"081B4A", x"000B2E", x"23395A", x"0A1C3A", x"BECED9", x"000126", x"F8FFF7", x"0A0C39", x"022245", x"021C43", x"3F4C6D", x"000223", x"061940", x"0C234A", x"031846", x"021E44", x"032341", x"021E4A", x"000820", x"FFFCFF", x"F8FFFF", x"36465B", x"E2F4F7", x"F4F9FA", x"FFFEFF", x"FBFEF7", x"F9FFF5", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFF9", x"1A2144", x"EEFFFF", x"FFFDE7", x"BBC6D5", x"00002E", x"022040", x"011A47", x"021E47", x"01163D", x"0A1F47", x"000A35", x"F0FFFF", x"040D37", x"091650", x"011835", x"FFFBFE", x"0B0D31", x"021340", x"FFF8FF", x"090021", x"011A4A", x"7D8DA0", x"303E65", x"021C41", x"000732", x"021549", x"05002E", x"0A1E49", x"022141", x"081C44", x"061C46", x"021D43", x"052340", x"0A174A", x"13203E", x"405F87", x"061239", x"42486E", x"273A5F", x"021D41", x"071540", x"071843", x"DFE0FC", x"0A1135", x"0A1C43", x"0A1C49", x"162851", x"909EB0", x"011540", x"022140", x"0B1646", x"041F45", x"091C43", x"0D1036", x"FAFFFE", x"FCFCFC", x"1E2A52", x"EEFAFB", x"FAFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFEFB", x"FCFDFA", x"40506F", x"BDBFDB", x"FAFBFF", x"FEFFFF", x"000029", x"022145", x"031E43", x"081E45", x"011B43", x"041F48", x"1B2046", x"7F839C", x"0B052F", x"4E627A", x"9999BA", x"0A1943", x"011746", x"D3DFEA", x"070F39", x"010127", x"8998AE", x"000F2F", x"090B2F", x"A9BAD6", x"232F4A", x"A2B3C8", x"2D3A52", x"0A214C", x"071D4A", x"021F43", x"011842", x"011A44", x"091A3D", x"F8FDFE", x"010B2F", x"022046", x"060330", x"8599AC", x"0C1B4B", x"021F43", x"041F4B", x"061335", x"EEF4F7", x"000C36", x"072144", x"0A1941", x"011842", x"021A43", x"0A1E49", x"081E4A", x"0A0931", x"475877", x"FFFEF9", x"FFFEF9", x"050B31", x"F0FFFF", x"FFFFFF", x"FFFDF9", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FEFFF5", x"FDFEF7", x"FDFFFB", x"9B9EBE", x"495468", x"FBFFFF", x"F6FFFC", x"363A5D", x"001138", x"081E4A", x"021F47", x"071C42", x"031C45", x"05052A", x"314579", x"0A0E40", x"091843", x"022043", x"021F44", x"7585A1", x"000A30", x"C3C6DB", x"01112B", x"000C2E", x"FEFEFF", x"04002D", x"0A194B", x"02103B", x"F7F9FF", x"00072D", x"081C42", x"031E44", x"072047", x"091B42", x"021B46", x"3E537A", x"3A5875", x"071D40", x"011A42", x"97A5B7", x"011336", x"021D44", x"071A49", x"13143B", x"C0C7E0", x"1D2F55", x"02214D", x"031B3C", x"021E3E", x"021F44", x"061E4B", x"000822", x"D4D6E5", x"F5FFFF", x"FEFEFE", x"000225", x"FEFFFC", x"FEFEFE", x"FEFFFF", x"FAFDFB", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FEFEFF", x"F6F8F0", x"FEFAF4", x"FAFCF4", x"FAFBFE", x"04092C", x"FFFEFB", x"FFFEFB", x"CFDBEA", x"00001D", x"071C43", x"0A1942", x"021F4A", x"081A49", x"021D4B", x"061E4B", x"081C46", x"0A214A", x"021D40", x"35496F", x"F9F5FE", x"00092B", x"031C40", x"000033", x"F8FFFA", x"0B113D", x"022042", x"011B46", x"A7B2AE", x"0F1F47", x"02213E", x"031F49", x"061B4C", x"021E42", x"081C44", x"010F35", x"EAF5F4", x"07123F", x"0B1539", x"838F9F", x"000B32", x"0A2048", x"022044", x"041F44", x"051743", x"0E1F48", x"051C43", x"031C45", x"031B44", x"000A32", x"303B59", x"FFFEFF", x"FAFBFF", x"A9B4BF", x"292E4F", x"FBFAFF", x"FEFBFF", x"FCFAFB", x"FFFFF9", x"FAFDF6", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FBFAF4", x"FAFAFC", x"232642", x"9DAFD4", x"FBFFFC", x"FBFFF4", x"696E8A", x"00052D", x"071D49", x"071D41", x"021E45", x"081C44", x"061A40", x"011944", x"011B41", x"163156", x"000F35", x"062045", x"081B43", x"01173D", x"F6FBFF", x"000017", x"011C47", x"000032", x"F2FFFF", x"010039", x"000D2E", x"021D4B", x"021D45", x"021D45", x"021D45", x"011C43", x"9FA3C1", x"CDCBD5", x"A0A5B1", x"232C4E", x"0C1D43", x"051B47", x"021D45", x"042042", x"071A4A", x"021E43", x"021C40", x"061340", x"0A102F", x"EAEDF6", x"FFFFF4", x"FFFCFE", x"141C39", x"C5C6DF", x"FEFEF4", x"FFFEFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"F4F4F4", x"FEFBFC", x"FBFFFC", x"D2DFE6", x"0A1231", x"FEFFFA", x"FBFEFC", x"FFFBFF", x"4B5A75", x"00002E", x"021C40", x"051B47", x"021E4A", x"021E46", x"021C42", x"091F49", x"091D45", x"032048", x"011B42", x"011C42", x"000030", x"B3B8D2", x"697CA1", x"92A6A8", x"0A0332", x"020A2D", x"F6FFFF", x"000038", x"021D45", x"021D45", x"021D45", x"031E46", x"011847", x"020027", x"000732", x"06214D", x"071E47", x"021F43", x"021E47", x"061E4B", x"022346", x"041137", x"070F3E", x"C8C6CE", x"FDFEFF", x"FCF7F6", x"838C9F", x"24294A", x"F8FFFF", x"FFFFFC", x"FCFAFE", x"FEFEFB", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FCFCFC", x"FFFFFC", x"FFFFFC", x"FEFEFF", x"FEFCFF", x"556377", x"2F3A60", x"F9FFFE", x"FFFBFF", x"FEFFF1", x"787F95", x"04052E", x"000E36", x"062141", x"021F44", x"07194B", x"021E46", x"021D45", x"091F49", x"0A1E4B", x"021D42", x"081C46", x"07173C", x"011C4D", x"021D42", x"0A1841", x"666997", x"0C113A", x"021D45", x"021D45", x"021D45", x"021D45", x"071F42", x"091E48", x"092346", x"022047", x"011A46", x"022041", x"0A1C42", x"00042F", x"1E2A51", x"EBE6E2", x"FAFDF9", x"FFFFFF", x"C7CEE2", x"0C1433", x"F3FFFF", x"FCFBFF", x"FFFFFF", x"FBFAF7", x"FBFBFB", x"FAFDFB", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FEFEFB", x"FFFFFC", x"FFFFFF", x"FFFFFC", x"FEF9F5", x"F8FFFA", x"FBF7FF", x"3B4C65", x"303A54", x"FAFFF9", x"FBFAFF", x"FBFFF6", x"F0EAFE", x"3C496D", x"000A2D", x"090E2F", x"0A1D45", x"061941", x"022044", x"011B40", x"031C41", x"051A40", x"021F44", x"0A1B4A", x"071E45", x"0A2054", x"01193B", x"03263F", x"021D45", x"021D45", x"021D45", x"021D45", x"021C46", x"022043", x"011841", x"02183E", x"000627", x"101B40", x"8895B0", x"FFFEFF", x"FFF7FF", x"F6FFFF", x"ACB6BE", x"0F1336", x"C8CEE2", x"F5FDF7", x"FFFDF9", x"F9FFFF", x"FFFCFE", x"FEFEFE", x"F9F9F6", x"FCFCFC", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"F9FFF6", x"6C7093", x"151C3C", x"ABBFDA", x"FFFEFF", x"FEFFFF", x"FEFEFE", x"FFFAFF", x"898FA8", x"1D3758", x"001037", x"010026", x"000C32", x"01163E", x"021D47", x"021C44", x"021D47", x"021D47", x"021E48", x"021D47", x"021E46", x"011A42", x"011139", x"000A2E", x"00002A", x"031940", x"435777", x"C8C2D7", x"FFFCFF", x"FBFEFC", x"FAFFFF", x"FFFFFF", x"4D5B75", x"171A3E", x"E2E5FB", x"FDFFEA", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFCFF", x"FEFFF9", x"F6F7FA", x"EBEDFC", x"283056", x"222952", x"ADBCC7", x"F3FFF7", x"FEFFFC", x"FFFAFF", x"FFFAFA", x"FFFEF6", x"FEFFFF", x"CAD6E1", x"96A8B4", x"798997", x"61778D", x"54687E", x"576C83", x"697F96", x"8396A4", x"A3B3BD", x"EBEEF7", x"FFF8FE", x"FFFDFA", x"FFF4FF", x"FFFCFF", x"FBFEF7", x"F3FFFF", x"56607D", x"11183E", x"687696", x"FBFEFF", x"FFFFFC", x"FBFAF5", x"FFFEFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFC", x"FAFCF4", x"FDFEF7", x"FFFFFF", x"FDFEFF", x"FAFAF7", x"F0FAFE", x"555F80", x"12234B", x"25385F", x"8094A7", x"DAE9E9", x"F8FFFA", x"FBFFFF", x"FBFBF9", x"FFFEFA", x"FEFFFA", x"FDFFF9", x"FEFFFA", x"FEFFFA", x"FAFDF6", x"FDFFFB", x"FEFFFC", x"FFFFFA", x"ADC2C7", x"4B5E7E", x"1A2A55", x"1B2C55", x"94A2B8", x"FBFFFC", x"FEFBFF", x"FFFFFC", x"FFFFFA", x"FBFDF5", x"FFFFFC", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FEFEFE", x"FFFFFF", x"FAFDFB", x"FEFFFF", x"FFFCFF", x"FBFFFF", x"FEFFFC", x"FFF8FF", x"FFFFF6", x"FFFEFA", x"F8FDFB", x"C1D4D0", x"6D7991", x"3A4C6B", x"1A3156", x"122C52", x"122B53", x"122B53", x"112A52", x"122B53", x"133053", x"243A5B", x"4C5874", x"8F93AD", x"E8F3EF", x"FFFEFC", x"FAF6F0", x"FDFFF2", x"FFFAFF", x"F9FEFC", x"FEFFFF", x"FFFEFC", x"FEFFFF", x"FCFCFC", x"FAFAFA", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", x"FFFFFF", 
x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"
);

	
begin

	-- Add user logic here
	int_X_Coord <= unsigned(X_Cord);
	int_Y_Coord <= unsigned(Y_Cord);
	int_X_Orig <= unsigned(slv_reg0);
    int_Y_Orig <= unsigned(slv_reg1);
    img_width <= unsigned(slv_reg2);
    img_height <= unsigned(slv_reg3);
	
	use_image <= '1' when int_X_Coord >= int_X_Orig and 
	                      int_X_Coord < int_X_Orig + img_width and
						  int_Y_Coord >= int_Y_Orig and 
						  int_Y_Coord < int_Y_Orig + img_height
				  else '0';
	
	image_next_index <= to_integer((int_Y_Coord-int_Y_Orig)*img_width + (int_X_Coord-int_X_Orig)) when use_image='1' else 0;
	image_next_pixel <= image(image_next_index);
	
	--rgb_next <= RGB_IN_I;
	
	rgb_next <= image_next_pixel when use_image = '1' else RGB_IN_I;
	RGB_IN_O 	<= rgb_next;
	
	VDE_IN_O	<= VDE_IN_I;
	HB_IN_O		<= HB_IN_I;
	VB_IN_O		<= VB_IN_I;
	HS_IN_O		<= HS_IN_I;
	VS_IN_O		<= VS_IN_I;
	ID_IN_O		<= ID_IN_I;
	
	slv_reg0out <= slv_reg0;
	slv_reg1out <= slv_reg1;
	slv_reg2out <= slv_reg2;
	slv_reg3out <= slv_reg3;
	slv_reg4out <= slv_reg4;
	slv_reg5out <= slv_reg5;
	slv_reg6out <= slv_reg6;
	slv_reg7out <= slv_reg7;

end Behavioral;